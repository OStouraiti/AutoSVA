bind riscv_CoreReorderBuffer riscv_CoreReorderBuffer_prop
	#(
		.ASSERT_INPUTS (0)
	) u_riscv_CoreReorderBuffer_sva(.*);