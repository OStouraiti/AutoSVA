bind imuldiv_IntMulDivIterative imuldiv_IntMulDivIterative_prop
	#(
		.ASSERT_INPUTS (0)
	) u_imuldiv_IntMulDivIterative_sva(.*);