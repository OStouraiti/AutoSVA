bind riscv_Core riscv_Core_prop
	#(
		.ASSERT_INPUTS (0)
	) u_riscv_Core_sva(.*);