bind imuldiv_IntDivIterative imuldiv_IntDivIterative_prop
	#(
		.ASSERT_INPUTS (0)
	) u_imuldiv_IntDivIterative_sva(.*);