bind imuldiv_IntMulIterative imuldiv_IntMulIterative_prop
	#(
		.ASSERT_INPUTS (0)
	) u_imuldiv_IntMulIterative_sva(.*);